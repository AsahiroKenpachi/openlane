module inverter (input a, output wire b);
not(b,a);
//assign b=~a;
endmodule
